.title KiCad schematic
.include "C:\Users\Elvis\3D Objects\Electronique\KICAD\KICAD 6\test_kicad_amelioration\54act00.lib"
.model mult_1 el_mult(in_offset =[0.1 0.1]
+ in_gain =[10.0 10.0] out_gain =5.0 out_offset =0.05)

V1 in1 GND pulse(0 5 2n 2n 2n 50u 100u)
V2 in2 GND sin(0 1 10k 30u)
a1 [in1 in2] Net-_R1-Pad1_ mult_1
R1 Net-_R1-Pad1_ GND 0.1
.save @v1[i]
.save @v2[i]
.save @r1[i]
.save V(Net-_R1-Pad1_)
.save V(in1)
.save V(in2)
.tran 1u 600u

.end

